module andgate(input [2:0] a,
           output y);

    assign y = &a;

endmodule