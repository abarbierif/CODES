module buffer(a, y);

    input a;
    output y;

    assign y = a;

endmodule

